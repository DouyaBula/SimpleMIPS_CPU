// baudrate = clk_freq / num_cycles
`define PERIOD_BAUD_9600    16'd2604    // PERIOD = 10^9ns / 9600baud / 40ns(25MHz)  
`define PERIOD_BAUD_38400   16'd651
`define PERIOD_BAUD_57600   16'd434
`define PERIOD_BAUD_115200  16'd217